`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/21/2021 08:19:09 PM
// Design Name: 
// Module Name: delay_counter_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module delay_counter_tb;

    logic clk, rst, delay_start, delay_done;
    
    delay_counter (.clk, .rst, .delay_start, .delay_done);
    
    
    
    

endmodule
